----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    12:50:00 03/13/2016 
-- Design Name: 
-- Module Name:    shift16 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity shift16 is
port(select_bit:in std_logic;
shift_type:in std_logic_vector(1 downto 0);
inp:in std_logic_vector(31 downto 0);
outp:out std_logic_vector(31 downto 0));
end shift16;

architecture Behavioral of shift16 is


begin

SHIFT:process(select_bit,inp)
begin
if (select_bit = '1') then
 case shift_type is
  when "00" =>
  --logic left
  outp(15 downto 0) <= "0000000000000000";
  outp(31 downto 16) <= inp(15 downto 0);
  when "01" =>
  --logic right
  outp(31 downto 16) <= "0000000000000000";
  outp(15 downto 0) <= inp(31 downto 16);
  when "11" =>
  --arith right
  outp(31) <= inp(31);
  outp(30) <= inp(31);
  outp(29) <= inp(31);
  outp(28) <= inp(31);
  outp(27) <= inp(31);
  outp(26) <= inp(31);
  outp(25) <= inp(31);
  outp(24) <= inp(31);
  outp(23) <= inp(31);
  outp(22) <= inp(31);
  outp(21) <= inp(31);
  outp(20) <= inp(31);
  outp(19) <= inp(31);
  outp(18) <= inp(31);
  outp(17) <= inp(31);
  outp(16) <= inp(31);
  outp(15 downto 0) <= inp(31 downto 16);
  when "10" =>
  outp(31 downto 16) <= inp(15 downto 0);
  outp(15 downto 0) <= inp(31 downto 16);
  when others =>
  outp <= inp;
 end case;
else
 outp <= inp;
end if;

end process;

end Behavioral;

